
module out_ram (
    input wire clk,
    input wire wen,             // ?????
    input wire [10:0] addr,      // ????
    input wire [11:0] data_in   // ????
);

    // ROM?????????784????8?
    reg [11:0] ram [0:1728];


    // ???
    always @(posedge clk) begin
        if (wen) begin
            ram[addr] <= data_in;  // ?ROM?????????????
        end
    end

endmodule

